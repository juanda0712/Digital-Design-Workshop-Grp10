module setting(output logic [5: 0] y);
	y = 1 & 1;
endmodule